`timescale 1ns/1ns
`include "mem_parameters.v"

module mem_tb ();